module sbox_combinational (x,sx);
 input[3:0] x;
 output reg [3:0] sx;
 always @(x)
 begin
 	sx= {(~x[3]&~x[1]& ~x[0]) | (~x[3]&x[1]&x[0]) | (~x[3]&x[2]&x[1]) | (x[3]&~x[2]&x[0]) | (x[3]&~x[2]&x[1]),
 	(~x[3]&~x[2]& ~x[1]) | (x[3]&x[2]&~x[1]) | (x[3]&~x[1]&x[0]) | (~x[2]&x[1]&~x[0]) | (~x[3]&x[2]&x[1]&x[0]),
 	(x[3]&~x[2]& ~x[1]) | (x[3]&x[2]&x[0]) | (~x[3]&~x[2]&x[1]) | (~x[3]&x[1]&~x[0]) | (~x[2]&x[1]& ~x[0]),
 	 (x[3]&x[1]& ~x[0]) | (~x[3]&~x[2]&x[0]) | (~x[3]&x[1]&x[0]) | (x[3]&~x[2]&~x[0]) | (~x[3]&x[2]& ~x[0] & ~x[1]) | (x[3]&x[2]& ~x[1] & x[0])};

 end
endmodule 